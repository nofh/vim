b0VIM 7.3      ���S�   �  dendev                                  lt-devos                                /mnt/awt/dev-denis/organisme/wp-content/plugins/wp_plugin_organisme/organisme.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �      M            
   N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ad  !   i     M   �  �  �  �  �  E  B  +    �  �  �  �  �  g  K  .  	  �  �  �  \  I  �  �  �  }    �  �  g  e    
  �
  l
   
  �	  �	  �	  c	  	  �  �  ?  &  �  q  e    �  �  �  V    �  �  ^    �  F  E  &  �  �  �  o  #  �  �  y  g  e    �  x  i  h                                   // renders 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/Import.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/CustomTinyMce.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/OrganismeAdmin.php'; { if( is_admin() )   *----------------------------------------------------------------------------*/  * ADMIN /*----------------------------------------------------------------------------* add_action( 'plugins_loaded', array( 'OrganismePublic', 'get_instance' ) ); // instancie le front  register_deactivation_hook( __FILE__, array( 'OrganismeCommun', 'deactivate' ) ); register_activation_hook( __FILE__, array( 'OrganismeCommun', 'activate' ) ); // activation et desactivation  require_once plugin_dir_path( __FILE__ ) . 'src/public/includes/shortcodes/OrganismesSHC.php'; require_once plugin_dir_path( __FILE__ ) . 'src/public/includes/shortcodes/OrganismeSHC.php'; require_once plugin_dir_path( __FILE__ ) . 'src/public/includes/shortcodes/ShortCode.php'; require_once plugin_dir_path( __FILE__ ) . 'src/public/OrganismePublic.php';  *----------------------------------------------------------------------------*/  * PUBLIC /*----------------------------------------------------------------------------* add_action( 'plugins_loaded', array( 'OrganismeCommun', 'get_instance' ) ); // instancie le commun   require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/taxos/TagTAXO.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/taxos/Taxonomie.php'; // taxonomy require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/OrganismeAPI.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/CustomPostTypeAPI.php'; // custom post types api require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/OrganismeCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/CustomPostType.php';  // custom post types require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/handlers/FormHandler.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/handlers/AjaxHandler.php'; // handlers // logeur -> require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/Db.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/Utils.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/OrganismeCommun.php';  *----------------------------------------------------------------------------*/  * COMMUN  /*----------------------------------------------------------------------------* }     require_once $emplacement_autoload; //require_once(): http:// wrapper is disabled in the server configuration by allow_url_include=0 { if( file_exists ( $emplacement_autoload ) ) $emplacement_autoload = plugin_dir_path( __FILE__ ) . 'src/commun/assets/vendor/autoload.php'; require_once plugin_dir_path( __FILE__ ) . 'src/config.php';  require_once plugin_dir_path( __FILE__ ) . 'src/config.php';  *----------------------------------------------------------------------------*/  * CONFIG & VENDOR /*----------------------------------------------------------------------------*   */  * Git Plugin URI: http://magneto/stash/projects/WPPLO/repos/wp_plugin_organisme/browse  * Text Domain:       organisme_lang  * Author:            dendev  * Version:           4.3.1  * Description:       Organismes ICT DigitalWallonia.be  * Plugin URI:        @TODO  * Plugin Name:       Organisme  * @wordpress-plugin  *  * @author   dendev <ddv@awt.be>  * @package  Structure  * @category Organisme  *  * also follow WordPress Coding Standards and PHP best practices.  * A foundation off of which to build well-documented WordPress plugins that  *  * WordPress Plugin Organisme. /** <?php ad  �  �     
   �  @  �  �  p      �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ?> }     add_action( 'plugins_loaded', array( 'OrganismeAdmin', 'get_instance' ) );      include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/OrganismeSAVE.php';     include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/CustomPostTypeSAVE.php';     // saves     include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/OrganismeRENDER.php';     include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/CustomPostTypeRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/AdminRENDER.php'; 