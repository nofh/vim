b0VIM 7.3      	��S�     dendev                                  lt-devos                                /mnt/awt/dev-denis/test/wp-content/plugins/wp_plugin_organisme/src/commun/includes/handlers/AjaxHandler.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �                  W               a                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ad  W  �        �  �  �  �  �  |  C    �  �  �  �  �  �  �  p  i  :  2    
  �  /  )  (        �  �  �  h  a  M  E      �  �  �  ~  u  \        �
  �
  �
  �
  e
  ^
  
  

  �	  �	  :	  3	  �  �  �  �  �  K    �  �  �  �  h  g  8    �  �  �  U  B    �  �  �  7  �  �    q  ^  0  �  �  �  y  K  �  �  M    �  �               case 'recuperer_valeurs_autocompletion': // pour bouton_generateurs.js             break;             $resultat['items'] = $db->recuperer_tags_deja_importer();         case 'recuperer_tags_deja_importer': // pour bouton_generateurs.js             break;             $resultat['items'] = $db->recuperer_cpt_localisations( $args['tag'], $args['post_type'], $args['post_id'], 'ASC', $args['certification_active'] );          case 'recuperer_infos_localisations':             break;             $resultat['totaux'] = $messages['totaux'];             $resultat['items'] = $messages['messages'];             $messages = $db->supprimer_cpts( $arg );         case 'supprimer_cpts': // pour import             break;             }                 $resultat['totaux'] = $messages['totaux'];                 $resultat['items'] = $messages['messages'];                 $messages = $db->ajouter_cpts( $cpts_importer );                 $cpts_importer = $import->importer_cpts_by_tag( $args['tag'], $args['limit'], $args['offset'], $message_import );                 $message_import = array();             {             if( is_array( $args ) )         case 'ajouter_cpts': // pour import             break;             $resultat['items'] = $import->recuperer_nb_cpts_a_importer( $arg ); // FIXME 1 represente rien         case 'recuperer_nb_cpts': // pour import         {         switch( $type_requete )         $resultat = array();         // choix de la rq devant etre executer          $import = new Import();         $db = Db::get_instance();         // init db          $args = ( ! empty( $_POST['args'] ) ) ? $_POST['args'] : false;         $arg = ( ! empty( $_POST['arg'] ) ) ? $_POST['arg'] : false;         $type_requete = str_replace( '_shortcode', '', $type_requete );         // formater args      {     private function executer_query( $type_requete )      */      * @return mixed[] le resultat avec ses infos completmentaires      *      * reformate le resultat en lui ajoutant le nb de resultat et la requete inital      * Choisi l'action adequate, sous traite le traitement       * Recupere les arguemnts de la demande, perapre le terrain      *      * @param $string type_requete le nom de la requete qui a etait demander      *      * Determine l'action a donner a une requete     /**      }        die( json_encode( $resultats, JSON_FORCE_OBJECT ) ); // FIXME nécessite version 5.3          // retourner l'info          $resultats = $this->executer_query( $type_requete );         // creer requete                  $type_requete = $_POST['type_requete'];          // recuperer l'info          global $wpdb; // this is how you get access to the database     {     public function executer_query_callback()       */      * @return null      *      * realise un die sur le resultat afin de l'envoyer a ajax      * et sous traite son traitement a executer_query      * recupere la demande       *      *  callback activer par wp     /**      }         add_action( 'wp_ajax_nopriv_executer_query', array( $this, 'executer_query_callback' ) ); // pour public          add_action( 'wp_ajax_executer_query', array( $this, 'executer_query_callback' ) ); // pour admin     {     public function __construct()      */      * Ajoute une action de recuperation ds wp      *      * Construct     /** { class AjaxHandle{ if{ if( ! class_exists( 'AjaxHandler' ) )   */  * les resultas renvoyer sont sous forme d'ojbect json  * renvoi le resultat plus la requete qui a etait demander a wp  * recup la demande et execute la fonction coorespondant  * Fonctionne pour la partie admin ou public  *  * Intercepete les requetes ajax faite a wp /** namespace Structure\Handlers; <?php ad  O  �        �  s    x  a  L        �  c  �  �  �  �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ?>???> }     }         }             return $resultat;             // fin              $resultat['requete'] = array( 'type_requete' => $type_requete, 'arg' => $arg, 'args' => $args );             $resultat['count'] = ( array_key_exists( 'items', $resultat ) ) ? count( $resultat['items'] ) : false;             // ajout des infos de la requete au resultat              }                 $resultat['items'] = 'vide';              default:                 break;                 $resultat['items'] = $db->recuperer_cpt_by_post_title_or_name_contact( $args['nom_champ'], $args['valeur_rechercher'], $args['post_type'] );             case 'recuperer_cpt_by_post_title_or_name_contact': // pour bouton_generateurs.js                 break;                 $resultat['items'] = $db->recuperer_valeurs_autocompletion( $args['nom_champ'], $args['post_type'] ); ad  _   �     W   �  �  �  �  �  �  y  S  I  �  f  \  [  O  +        �  �  x  `  T  !    �  �  �  y  x  [      �  �  �  �  �  K  @  �
  �
  �
  `
  
  �	  �	  �	  q	  g	  I	  �  �  h  g  P  *      �  �  �    J  �  �  �  l  Z  +  �  `     �  �  �  �  M    �  �  �  �  �  �  9  "  �                                                                                                             case 'recuperer_valeurs_autocompletion': // pour bouton_generateurs.js                 break;                 $resultat['items'] = $db->recuperer_tags_deja_importer();             case 'recuperer_tags_deja_importer': // pour bouton_generateurs.js                 break;                 $resultat['items'] = $db->recuperer_cpt_localisations( $args['tag'], $args['post_type'], $args['post_id'], 'ASC', $args['certification_active'] );              case 'recuperer_infos_localisations':                 break;                 $resultat['totaux'] = $messages['totaux'];                 $resultat['items'] = $messages['messages'];                 $messages = $db->supprimer_cpts( $arg );             case 'supprimer_cpts': // pour import                 break;                 }                     $resultat['totaux'] = $messages['totaux'];                     $resultat['items'] = $messages['messages'];                     $messages = $db->ajouter_cpts( $cpts_importer );                     $cpts_importer = $import->importer_cpts_by_tag( $args['tag'], $args['limit'], $args['offset'], $message_import );                     $message_import = array();                 {                 if( is_array( $args ) )             case 'ajouter_cpts': // pour import                 break;                 $resultat['items'] = $import->recuperer_nb_cpts_a_importer( $arg ); // FIXME 1 represente rien             case 'recuperer_nb_cpts': // pour import             {             switch( $type_requete )             $resultat = array();             // choix de la rq devant etre executer              $import = new Import();             $db = Db::get_instance();             // init db              $args = ( ! empty( $_POST['args'] ) ) ? $_POST['args'] : false;             $arg = ( ! empty( $_POST['arg'] ) ) ? $_POST['arg'] : false;             $type_requete = str_replace( '_shortcode', '', $type_requete );             // formater args          {         private function executer_query( $type_requete )          */          * @return mixed[] le resultat avec ses infos completmentaires          *          * reformate le resultat en lui ajoutant le nb de resultat et la requete inital          * Choisi l'action adequate, sous traite le traitement           * Recupere les arguemnts de la demande, perapre le terrain          *          * @param $string type_requete le nom de la requete qui a etait demander          *          * Determine l'action a donner a une requete         /**          }             die( json_encode( $resultats, JSON_FORCE_OBJECT ) ); // FIXME nécessite version 5.3              // retourner l'info              $resultats = $this->executer_query( $type_requete );             // creer requete              $type_requete = $_POST['type_requete'];              // recuperer l'info              global $wpdb; // this is how you get access to the database         {         public function executer_query_callback()           */          * @return null          *          * realise un die sur le resultat afin de l'envoyer a ajax          * et sous traite son traitement a executer_query          * recupere la demande           *          *  callback activer par wp         /**          }             add_action( 'wp_ajax_nopriv_executer_query', array( $this, 'executer_query_callback' ) ); // pour public              add_action( 'wp_ajax_executer_query', array( $this, 'executer_query_callback' ) ); // pour admin         {         public function __construct()          */          * Ajoute une action de recuperation ds wp          *          * Construct         /**     {     class AjaxHandler 