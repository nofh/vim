b0VIM 7.3      z(�S;�   dendev                                  lt-devos                                ~dendev/public_html/NeaLoca/wp-content/plugins/fmwp/src/config.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �      /                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ad  �	  �
     /   �  �  �  �  �  �  �  �  �  ~  `  ?  >  4  �  �  �  �  o  H  G  9        �    2  �  �  �  �  G    �  �  �  w  4  3  )  (      �
  �
  �
  �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ???> error_reporting(E_ALL); define('WP_DEBUG_LOG', true); define('WP_DEBUG', true); // debug  // global  define( 'EMP_VENDORS', URL_PLUGIN . 'src/commun/assets/vendors/'); // vendors  define( 'EMP_IMG_ADMIN', URL_PLUGIN . 'src/admin/assets/img/'); define( 'EMP_IMG_PUBLIC', URL_PLUGIN . 'src/public/assets/img/'); define( 'EMP_IMG_PUBLIC', URL_PLUGIN . 'src/commun/assets/img/'); define( 'URL_PLUGIN', plugins_url() . '/fmwp/'); // FIXME define( 'URL_PLUGIN', plugins_url() . '/' . dirname( plugin_basename( __FILE__ ) ) . '/' ); // Img    define( 'EMP_ADMIN_VIEWS', plugin_dir_path( __FILE__ ) . 'admin/views/' ); define( 'EMP_PUBLIC_VIEWS', plugin_dir_path( __FILE__ ) . 'public/views/' ); define( 'EMP_COMMUN_VIEWS', plugin_dir_path( __FILE__ ) . 'commun/views/' ); define( 'EMP_PLUGIN', plugin_dir_path( __FILE__ ) ); // emplacement  define( 'TEXT_DOMAIN', 'fmwp_langue' ); // traduction  define( 'TAXO_LANGUE', 'LangueTaxo' ); define( 'TAXO_TEST', 'TestTaxo' ); // Taxonomie  define( 'PREFIX_META', '_fw_' ); // TODO passer de _ec vers og define( 'PREFIX_PLUGIN', 'fw_' ); // TODO readapation voir creation cpt pour le nom  // prefix  define( 'PLUGIN_SLUG', 'fmwp' ); define( 'VERSION', '1.0.0' ); // Version   */  * @author   dendev <ddv@awt.be>  * @package  Organisme  * @category Fmwp  *  * Configuration du plugin /** <?php 