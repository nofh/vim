b0VIM 7.3      K��S�5  =G  dendev                                  lt-devos                                /mnt/awt/dev-denis/test/wp-content/plugins/wp_plugin_organisme/src/commun/includes/Utils.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �      l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ad  �  Y     l   �  �  �  �  �  �  �  v  l  L  >  �  �  �  �  �  r  g    �  �  �  �  N  B    �  �  �  �  l  ^      �  �  �  �  �  �  �  Q  G  *  )    �
  �
  �
  �
  f
  T
  
  	
  �	  �	  �	  �	  �	  s	  a	  F	  4	  &	  %	  		  �  �  �  �  �  �  w  L  K      �  �  �  �  M  .        �  �  �  �  �  �  y  o  n  &         �  �  �  �  �  k  a  [  Y  X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   }     }         }             return $etic;              }                 $etic = true;             {             if( $nom_tag == 'charte_etic' || $nom_tag == '24' )              $etic = false;         {         public static function is_tag_etic( $nom_tag ) // @depreacted ?          }             return $slug_tag;              }                 }                     break;                 {                 if( $slug_tag )                  }                     }                         break;                         $slug_tag = $tag->message;                     {                     if( $tag->id_tag == $id_tag )                 {                 foreach( $tags_categorie as $tag )             {             foreach( $tags as $tags_categorie )              $tags = $db->recuperer_tags();             $db = Db::get_instance();              $slug_tag = false;         {         public static function get_slug_tag( $id_tag )          }             return $id_tag;              }                 }                     break;                 {                 if( $id_tag )                  }                     }                         break;                         $id_tag = $tag->id_tag;                     {                     if( $tag->message == $slug_tag )                 {                 foreach( $tags_categorie as $tag )             {             foreach( $tags as $tags_categorie )              $tags = $db->recuperer_tags();             $db = Db::get_instance();              $id_tag = false;         {         public static function get_id_tag( $slug_tag )          }             return $ids_cpt_sticky;              }                 }                      $ids_cpt_sticky[] = $id_sticky;                 {                 if( get_post_type( $id_sticky ) === $nom_cpt )             {             foreach( $ids_sticky as $id_sticky )             $ids_cpt_sticky = array();              $ids_sticky = get_option( 'sticky_posts' );         {         public static function get_sticky_cpts( $nom_cpt )          */          * @return string[] contenant les ids des custom post types sticky          *          * @params string $nom le nom du custom post type ( ex: organisme );          *          * et etant sticky          * recupere les custom post type ayant pour nom la valeur passer en arg          *          * recupere les cpts sticky.         /**          }             }                 echo("<script>console.log('PHP: ".json_encode( print_r( $data ), JSON_HEX_APOS | JSON_HEX_QUOT )."');</script>");             {             if( self::$_debug )         {         public static function debug( $data )     {     class Utils { if( ! class_exists( 'Utils' ) )   namespace Structure\Commun; <?php 