b0VIM 7.3      jP�S�  �,  dendev                                  lt-devos                                /mnt/awt/dev-denis/organisme/wp-content/plugins/wp_plugin_organisme/src/commun/includes/Db.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp	 �      n         
   g   o         <   �         6           h   H        $   �        =   �     	   j           D   {                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ad     �     n   �  �  �  �  �  6  �  �  �  �  �  �  �  �  �  �  �  J  B        �  �  �  �  �  �  `  X  .  (     �  �  �  �  �  �  �      �  g  f  ;  #    �
  �
  �
  �
  ^
  H
  �	  �	  k	  j	  	  �  �  �  u  3    �  �  �  H  !  �  �  z  U    �  �  �  �  X  >  (      �  �  �  �  �  �  �  c  b  [  Z  �  �  �  �  ^  8    �  �  �  s  O  +    �  �                                'child_of'      => 0,              'hierarchical'  => true,              'parent'         => '',             'slug'          => '',              'fields'        => 'all',              'number'        => '',              'include'       => array(),             'exclude_tree'  => array(),              'exclude'       => array(),              'hide_empty'    => true,              'order'         => 'ASC',             'orderby'       => 'name',          $args = array(     {     public function recuperer_tags_deja_importer( $associatif=true ) // un tag qui existe et un tag ayant des organisme ( qui a etait importer )      }           return $tags_recuperer;           }             echo "erreur imposible de deserialiser le contenu de l'option"; // TODO log         {         else         }             }                 }                     }                         }                             $tags_recuperer['autres'][] = $tag_tmp;                          {                         else                         }                             }                                 $tags_recuperer['autres'][] = $tag_tmp;                              default:                                 break;                                 $tags_recuperer['appartenance'][] = $tag_tmp;                              case 'appartenance':                                 break;                                 $tags_recuperer['affiliation'][] = $tag_tmp;                              case 'affiliation':                             {                             switch( $tag_tmp->type )                         {                         if( property_exists( $tag_tmp, 'type' ) )                         // conserve l'object ds sa categorie                           $tag_tmp->checked = $checked;                         $tag_tmp->existe = $existe;                         // enrichie l object avec les informations deduites                          $checked = ( $existe ) ? 'checked' : '';                         $existe = ( $existe == null ) ? false : true;                         $existe = get_term_by( 'slug', $tag_tmp->message, TAXO_TAG );                     {                     if( property_exists( $tag_tmp, 'message' ) )                 {                  if( is_object( $tag_tmp ) )             {             foreach( $tags_tmp as $tag_tmp )         {         if( $tags_tmp )         // si la unserialisation a reussit          $tags_tmp = get_option( PREFIX_META . 'tags_cpts', false );         $tags_recuperer = array( 'appartenance' => array(), 'affiliation' => array(), 'autres' => array() );     {     static function recuperer_tags() // FIXME via tag name plutot que slug non ? le slug peut changer le nom pas      // recuperer     } 		return self::$_instance;          }             self::$_instance = new self;         {         if( self::$_instance == null )      {     public static function get_instance()      */      * @return int une instance sur la class ( pas vraiment un int ... )      *      * Implemente le patterns singleton     /**      }         $this->_db = $wpdb;         global $wpdb;     {     private function __construct()      */      * recupere le wpdb global et wp et se le met en attribut      *       * Construct encore et tj     /**       private $_db;     private static $_instance = null; { class Db  */  * classe singletion, s'intacie via Db::get_instance()  * Exception pour CustomPostTypeApi ( est ses descedants ) qui benefici d'un privilige d'autonomie  * Tout elements accedant a la db viens chercher ses infos ici  *  * Centralise les acces db /** <?php ad  !  E     D   �  �  }  |  N    �  �  �  �  �  �         �  �  �  �  �  6  0  �  �  �  �  �  f  e  )  (  '        �
  �
  �
  �
  p
  J
  @
  
  
  �	  �	  �	  �	  q	  c	  Y	  X	  D	  >	  =	  	  �  �  �  �  �  f  e  d  P  J  H  E  D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ?> }     }         return $ok;           $ok = ( is_object( $rez ) || ! $rez ) ? false : true;          $rez = wp_set_post_terms( $post_id, $tag, TAXO_TAG, true );          $ok = false;     {     private function _ajouter_tag_cpt( $tag, $post_id )      }         return $ok;          }             }                 }                     break;                     $ok = true;                 {                 if( $post_tag->slug == $slug_tag )             {             foreach( $post_tags as $post_tag )         {         if( count( $post_tags ) > 0 )         $post_tags = wp_get_post_terms( $post_id, TAXO_TAG );          $ok = false;     {     private function _cpt_possede_tag( $slug_tag, $post_id )      }         return $post_id;           $post_id = ( $post_id == null ) ? false : $post_id;          $post_id = $this->_db->get_var( $this->_db->prepare( "SELECT pm.post_id FROM " . $this->_db->postmeta . " pm INNER JOIN " . $this->_db->posts . " p ON p.ID = pm.post_id WHERE pm.meta_key = '%s' AND pm.meta_value = '%s' AND p.post_status = '%s' ", PREFIX_META . $meta_key, $meta_value, 'publish' ) );     {     private function _cpt_possede_meta( $meta_key, $meta_value )      }         return $this->_cpt_possede_meta( 'id_' . $post_type, $id_cpt );     {     private function _cpt_existe_en_db( $id_cpt, $post_type ) // TOD id_organisme, id_evenement ,....      // --      }         $this->_db->delete( $this->_db->posts, array( 'post_type' => 'organisme' ) );          // post organisme          $this->_db->query( "DELETE FROM " . $this->_db->postmeta . " WHERE meta_key LIKE '_og%' " );          // meta datas                   }             wp_delete_term( $term->term_id, TAXO_TAG );         {         foreach( $terms as $term )         $terms = get_terms( TAXO_TAG, 'orderby=count' );         // supprimer les terms de la taxonomi          }             delete_option( PREFIX_META . 'tags_autres' );             delete_option( PREFIX_META . 'tags_affiliation' ); ad  �	  z
     $   �  ~    �  �  �  �  �  q  c    �  �  �  ~  t  s  >  h  g  X  	    �  �  �  �  �  �  �  �  Z  Y    �
  z
  
  Q
  
  �	  �	  o	  n	  P	  8	  	  �  �  �  `  5  �  �  �  �  �  D  9  �  �  �  �  �  �  /           �  �  �  �  �  �  �  W  M  �  �      �  �  �  �  �  �  �  �  �  �  �  �  �  �  �      // formater      }                  return $colonne;           //$this->debug();         }             $colonne = $this->_db->get_col( $this->_db->prepare( "SELECT DISTINCT meta_value FROM ". $this->_db->postmeta ." WHERE meta_key = '%s' ORDER BY meta_value DESC", PREFIX_META . $nom_champ ) );         {            else         }             $colonne = $this->_db->get_col( $this->_db->prepare( "SELECT DISTINCT meta_value FROM ". $this->_db->postmeta ." WHERE meta_key = '%s' ORDER BY meta_value DESC", PREFIX_META . $nom_champ ) );             $nom_champ = 'nom_contact'; // pour fair semblant d'etre generic .... // FIXME         {         else if( $nom_champ == 'nom_prenom_contact' ) // !!!! CAS particulier nom  contact ds agenda == nom prenom         }             $colonne = $this->_db->get_col( $this->_db->prepare( "SELECT DISTINCT post_title FROM ". $this->_db->posts ." WHERE post_type = '%s'  ORDER BY post_title", $post_type ) );         {         if( $nom_champ == 'post_title' )          $colonne = array();     {     public function recuperer_valeurs_autocompletion( $nom_champ, $post_type )      }          return $post_id;            }              }                  update_post_meta( $post_id, PREFIX_META . $nom, $valeur ); // meta_key unique              {              else               }                  // rien car setter ds le post              {              if( $nom == 'titre' || $nom == 'description' )          {          foreach( get_object_vars( $cpt ) as $nom => $valeur )            $post_id = wp_insert_post($post);          // save en db          );              'post_type'  => $post_type // FIXME stupide !! on va recuper le post type comment ?               'post_title' => $post_title,               'post_status' => 'publish',               'post_content' => $post_content,              'post_date' => date( 'Y-m-d H:i:s' ),              'post_author' => 1,              'comment_status' =>  'closed',          $post = array(          // creation du post           unset( $cpt->$attribut_post_content );         $post_content = $cpt->$attribut_post_content;         $attribut_post_content = 'description_' . $post_type;               $post_title = (property_exists( $cpt, $attribut_post_title ) ) ? $cpt->$attribut_post_titl        $post_title = ( property_exists( $cpt, $attribut_post_title ) ) ? $cpt->$attribut_post_title : '';         $attribut_post_title = 'nom_' . $post_type;         // recuperation du titre a utiliser pout le post title           $post_type = $cpt->post_type;         // recup du post_type          $post_id = false;     {     public function ajouter_cpt( $cpt )      }         return $messages;          $messages = array('messages' => $tmp_messages, 'totaux' => $totaux ) ;         // fin          $totaux = array( 'nb_deja_existant' => $nb_deja_existant, 'nb_mis_a_jour' => $nb_mis_a_jour, 'nb_sauvegarder' => $nb_sauvegarder, 'nb_supprimer' => 0, 'nb_tags_supprimer' => 0, 'nb_erreur' => $nb_erreur );         // totaux des orgs ajouter, mis a jour, ....          }             $tmp_messages[] = $cpt_message;             }                 $nb_erreur++;                 $cpt_message['erreur'] = 1;                 $cpt_message['message'] = __( 'Echec: ajout de ', TEXT_DOMAIN ) . $post_title ;              {             if( ! $post_id )             // gestion des erreurs              }                 $nb_sauvegarder++;                 $cpt_message['sauvegarder'] = 1;                 $cpt_message['message'] =  $post_title . __( " création et ajout du tag", TEXT_DOMAIN );                 $post_id = $this->_ajouter_tag_cpt( $slug_tag, $post_id );                 $post_id = $this->ajouter_cpt( $cpt ); ad  �  �     =   �  �  �  U  �  �  �  �  ~  R  1  �  �  �  {      �  �  �  �    C  4    �  �  �  u  f  [  Z  Y  ?  9  8  �
  �
  �
  �
  �
  �
  �	  �	  ^	  T	  �  -  #    	  =  3        �  �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  // formater      }                  return $colonn    // formater      }                  return $colonne;           //$this->debug();         }             $colonne = $this->_db->get_col( $this->_db->prepare( "SELECT DISTINCT meta_value FROM ". $this->_db->postmeta ." WHERE meta_key = '%s' ORDER BY meta_value DESC", PREFIX_META . $nom_champ ) );         {            else         }             $colonne = $this->_db->get_col( $this->_db->prepare( "SELECT DISTINCT meta_value FROM ". $this->_db->postmeta ." WHERE meta_key = '%s' ORDER BY meta_value DESC", PREFIX_META . $nom_champ ) );             $nom_champ = 'nom_contact'; // pour fair semblant d'etre generic .... // FIXME         {         else if( $nom_champ == 'nom_prenom_contact' ) // !!!! CAS particulier nom  contact ds agenda == nom prenom         }             $colonne = $this->_db->get_col( $this->_db->prepare( "SELECT DISTINCT post_title FROM ". $this->_db->posts ." WHERE post_type = '%s'  ORDER BY post_title", $post_type ) );         {         if( $nom_champ == 'post_title' )          $colonne = array();     {     public function recuperer_valeurs_autocompletion( $nom_champ, $post_type )      }          return $post_id;            }              }                  update_post_meta( $post_id, PREFIX_META . $nom, $valeur ); // meta_key unique              {              else               }                  // rien car setter ds le post              {              if( $nom == 'titre' || $nom == 'description' )          {          foreach( get_object_vars( $cpt ) as $nom => $valeur )            $post_id = wp_insert_post($post);          // save en db          );              'post_type'  => $post_type // FIXME stupide !! on va recuper le post type comment ?               'post_title' => $post_title,               'post_status' => 'publish',               'post_content' => $post_content,              'post_date' => date( 'Y-m-d H:i:s' ),              'post_author' => 1,              'comment_status' =>  'closed',          $post = array(          // creation du post           unset( $cpt->$attribut_post_content );         $post_content = ( property_exists( $cpt, $attribut_post_content ) ) ? $cpt->$attribut_post_content : '';         $attribut_post_content = 'description_' . $post_type;         // recuperer le 2 elements pour l'utiliser comme titre          unset( $cpt->$attribut_post_title ); ad  %   �     h   �  �  �  �  �  �  �  �  �  Z  T  :  9  �  �  s  m  l  ]  3  -    }  |  h  4  3  !  �  �  �  �  �  �  l  P  3      �  �  �  �  �  �  _  ^    �
  �
  �
  k
  ]
  \
  
  �	  �	  �	  l	  ^	  ]	  *	  	  �  �  �  �  y  b  �  �  �  n  A    �  �  �  @  %      �  �  �  A  /  �  �  K  "    �  �  �  :  �  v  Q  ?  1       �  �                                                   // si eixte pas alors on le cree en db               {             else             }                 }                    $nb_mis_a_jour++;                    $cpt_message['mis_a_jour'] = 1;                    $cpt_message['message'] = $post_title . __( " existe deja en db mais avec un autre tag, ajout du nouveau tag", TEXT_DOMAIN );                    $post_id = $this->_ajouter_tag_cpt( $slug_tag, $post_id );                    // si existe mais pas mm tag alors ajoute a l'existant le tag de l'cpt en arg                 {                 else                 }                     $nb_deja_existant++;                     $cpt_message['deja_existant'] = 1;                     $cpt_message['message'] = $post_title . __( " existe deja en db avec le même tag", TEXT_DOMAIN );                     // si existe et mm tag alors rien                 {                 if( $this->_cpt_possede_tag( $slug_tag, $post_id ) )                 // si existe test si possede le mm tag que l'cpt en arg                  $cpt_message['post_id'] = $post_id;                 //              {             if( $post_id )             $post_id = $this->_cpt_existe_en_db( $id_cpt, $post_type ); // id_cpt est l'id de organisme, id de evenemnt ...             // test si cpt existe deja en db              $cpt_message['erreur'] = -1;             $cpt_message['sauvegarder'] = -1;             $cpt_message['mis_a_jour'] = -1;             $cpt_message['deja_existant'] = -1;             // etat d'un cpt              $cpt_message = array( 'id' => $id_cpt, 'nom' => $post_title, 'message' => '', 'tag' => $slug_tag );//FIXME id devrait s'appeler id_cpt ( depend de 'api )             // message                          }                 $id_cpt = $cpt->$attribut_id_cpt;             {             if( property_exists( $cpt, $attribut_id_cpt ) )             $id_cpt = '';             $attribut_id_cpt = 'id_' . $post_type;              }                 $post_content = $cpt->$attribut_post_content;             {             if( property_exists( $cpt, $attribut_post_content ) )             $post_content = '';             $attribut_post_content = 'description_' . $post_type;              }                 $post_title = $cpt->$attribut_post_title;             {             if( property_exists( $cpt, $attribut_post_title ) )             $post_title = '';             $attribut_post_title = 'nom_' . $post_type; // FIXME pas generic              $post_type = $cpt->post_type;             // infos de base du post          {         foreach( $cpts as $cpt )          $tmp_messages = array();          // tout les messages          $nb_erreur = 0;         $nb_sauvegarder = 0;         $nb_mis_a_jour = 0;         $nb_deja_existant = 0;         // totaux     {     public function ajouter_cpts( $cpts, $slug_tag)      }         add_option( PREFIX_META . 'tags_cpts', $tags, '', false );         //ajouter          delete_option( PREFIX_META . 'tags_cpts' );         // nettoyer          $tags_formater = $this->formater_tags( $tags, true ); // TODO pas util car resultat simple ( a priori ) a fixer quand le webservice envera les tags         // formater     {     public function ajouter_tags( $tags )     // ajouter      }         return $post_id;          $post_id = $this->_db->get_var( $this->_db->prepare( "SELECT ID FROM " . $this->_db->posts . " WHERE post_title = '%s' AND post_type = '%s'", $nom, $post_type ) );          $post_id = false;     {     public function recuperer_id_par_post_title( $nom, $post_type )      }         return $ids;           //$this->debug();         }             }                 } ad  	   �      6   j    �  Q  �  �  [  E  ,    �  �  %  �  �  J    �
  t
  
  �	  �	  �	  �	  �	  L	  6	  �  �  �  D    �  =  �  U  �  �  V    �  c  M  4  �  E  �  �  6  �  �  �    �   �                            }                             . "ORDER BY pm.meta_value $ordre_trie", $post_type, $id_tag->term_taxonomy_id, $clee_trie ) );                             . "AND pm.meta_key ='%s' "                             . "AND r.term_taxonomy_id = '%s' "                             . "WHERE p.post_type = '%s' "                             . "INNER JOIN " . $this->_db->postmeta . " pm ON pm.post_id = p.id "                             . "INNER JOIN " . $this->_db->posts . " p ON p.id = r.object_id "                             . "FROM  " . $this->_db->term_relationships . " r "                         $ids = $this->_db->get_col( $this->_db->prepare( "SELECT p.id AS post_id, p.post_title AS post_title, pm.meta_key AS meta_key, pm.meta_value AS meta_value "                     { // etic avec certif autre que toute                     else                     }                            $certification_active,  $clee_trie, $id_tag->term_taxonomy_id, $post_type, $ordre_trie ) );                             "ORDER BY pmm.meta_value $ordre_trie ",                             "AND p.post_type = '%s' " .                             "WHERE tr.term_taxonomy_id = '%s' " .                             "INNER JOIN wp_terms ts ON ts.term_id = t.term_id " .                             "INNER JOIN wp_term_taxonomy t ON t.term_taxonomy_id = tr.term_taxonomy_id " .                             "INNER JOIN wp_term_relationships tr ON tr.object_id = p.id " .                             "INNER JOIN ( SELECT post_id, meta_value FROM wp_postmeta WHERE meta_key = '%s' ) pmm ON pmm.post_id = p.ID " .                             "INNER JOIN ( SELECT post_id, meta_value FROM wp_postmeta WHERE meta_key = '%s'  AND meta_value = '1' ) pm ON pm.post_id = p.ID " .                             "FROM wp_posts p " .                             "SELECT DISTINCT p.id " .                         $ids = $this->_db->get_col( $this->_db->prepare(                           // clee de trie est recut avec deja PREFIX_META                         $certification_active = PREFIX_META . $certification_active . '_etic';                     {                     if( $certification_active != 'toute' )                 {                 else // pour le trie sur les champs non post_title et non date                  }                      }                             . "ORDER BY STR_TO_DATE(  pm.meta_value, '%d.%m.%Y' ) $ordre_trie" );                             . "AND pm.meta_key = '${clee_trie}' "                             . "AND r.term_taxonomy_id = '${term_taxonomy_id}' "                             . "WHERE p.post_type = '${post_type}' "                             . "INNER JOIN wp_postmeta pm ON pm.post_id = p.id "                             . "INNER JOIN wp_posts p ON p.id = r.object_id "                             . "FROM wp_term_relationships r "                         $ids = $this->_db->get_col( "SELECT id, IFNULL( pm.meta_key, '00.00.0000' ) "                         $term_taxonomy_id = $id_tag->term_taxonomy_id;                         // etic( toute ) ou pas avec trie sur date                     {                      else                     }                             "ORDER BY STR_TO_DATE( pmm.meta_value, '%d.%m.%Y' ) $ordre_trie " );                             "AND p.post_type = '${post_type}' " .                             "WHERE tr.term_taxonomy_id = '${term_taxonomy_id}' " .                             "INNER JOIN wp_terms ts ON ts.term_id = t.term_id " .                             "INNER JOIN wp_term_taxonomy t ON t.term_taxonomy_id = tr.term_taxonomy_id " .                             "INNER JOIN wp_term_relationships tr ON tr.object_id = p.id " .                             "INNER JOIN ( SELECT post_id, meta_value FROM wp_postmeta WHERE meta_key = '${clee_trie}' ) pmm ON pmm.post_id = p.ID " . ad  2   6     <   �  �  �  �  �  N  M  5  4  �  �  �  �  f  X  W  �  �      �  �  <    ^
  
  �	  E	  	  �  F  0      �  2  �  �  [  �  �  �  :  (  �  _  #    �  �  �  n  V    �  �  j    �  6  5                                                                            "INNER JOIN ( SELECT post_id, meta_value FROM wp_postmeta WHERE meta_key = '${certification_active}'  AND meta_value = '1' ) pm ON pm.post_id = p.ID " .                             "FROM wp_posts p " .                         $ids = $this->_db->get_col( "SELECT DISTINCT p.id " .                         $term_taxonomy_id = $id_tag->term_taxonomy_id;                          $certification_active = PREFIX_META . $certification_active . '_etic';                         // etic avec certif active et trie sur date                      {                       if( $certification_active != 'toute' )                      }                         $clee_trie = PREFIX_META . 'date_souscription_etic';                     {                     if( $slug_tag == CHARTE_ETIC_TAG_NAME )                     $clee_trie = PREFIX_META . 'date_creation_organisme';                     // choix de la date selon est etic ou pas ( etic fonction avec souscription, non etic avec date creation )                 {                 else if( str_replace( PREFIX_META, '', $clee_trie ) == 'date_creation_ou_souscription_etic' ) // trie sur les champs dates                 }                     }                             . "ORDER BY p.post_title $ordre_trie", $post_type, $id_tag->term_taxonomy_id ) );                             . "AND r.term_taxonomy_id = '%s' "                             . "WHERE p.post_type = '%s' "                             . "INNER JOIN " . $this->_db->posts . " p ON p.id = r.object_id "                             . "FROM  " . $this->_db->term_relationships . " r "                         $ids = $this->_db->get_col( $this->_db->prepare( "SELECT p.id AS post_id, p.post_title AS post_title "                     {                     else                     }                             . "ORDER BY p.post_title $ordre_trie", $certification_active, $id_tag->term_taxonomy_id, $post_type ) );                             . "AND p.post_type = '%s' "                             . "WHERE tr.term_taxonomy_id = '%s' "                             . "INNER JOIN wp_terms ts ON ts.term_id = t.term_id "                             . "INNER JOIN wp_term_taxonomy t ON t.term_taxonomy_id = tr.term_taxonomy_id "                             . "INNER JOIN wp_term_relationships tr ON tr.object_id = p.id "                             . "INNER JOIN ( SELECT post_id, meta_value FROM wp_postmeta WHERE meta_key = '%s'  AND meta_value = '1' ) pm ON pm.post_id = p.ID  "                                         . "FROM wp_posts p "                         $ids = $this->_db->get_col( $this->_db->prepare( "SELECT DISTINCT p.id AS post_id "                          $certification_active = PREFIX_META . $certification_active . '_etic';                     {                     if( $certification_active != 'toute' ) // les non etic sont a certification_active == toute par defaut ( et mm par obligation voir bridage ds le shortcode organismes )                 {                 if( str_replace( PREFIX_META, '', $clee_trie ) == 'post_title' ) // trie sur le post_title              {             if( property_exists( $id_tag, 'term_taxonomy_id' ) )         {         if( is_object( $id_tag ) )          $id_tag = get_term_by( 'name', $slug_tag, TAXO_TAG );//Utils::get_id_tag( $slug_tag );          $ids = array();          $clee_trie = ( ! strstr( PREFIX_META, $clee_trie ) ) ? PREFIX_META . $clee_trie : $clee_trie;     {     public function recuperer_posts_ids_cpt( $slug_tag, $post_type, $clee_trie, $ordre_trie = 'ASC', $type_trie = 'string', $certification_active = 'toute' ) //TODO pas d'appel direct -> wp_post mais passer par db->post      */      *      * @return string[] ids renvoi tout les post_id des custom post type cpt selectionner  ad  +   �     j   �  �  �  {  z  Y  O  �  �  >  =  �  �  �  �  �  �  i  2  $  �  �  �  j  `  _  @  :  9  -      �  �  �  �  �  �  Y      �
  �
  �
  �
  �
  �
  �
  _
  ^
  &
  �	  �	  �	  �	  �	  �	  R	  %	  	  �  T  S  .  �  �  s  O  �  �  �  E  D  �  �  �  w  b  P  �  �  |  j  i  A  3  )      �  �  z  V  L  �  �  �  �  �  �  f  `  E  1  '  �  �                                                     delete_option( PREFIX_META . 'tags_appartenance' );         {         if( $tags )         // supprimer tags      {     public function supprimer_tout($tags=false)      }         return array( 'messages' => $messages, 'totaux' => $totaux );           $totaux = array( 'nb_supprimer' => $nb_supprimer, 'nb_tags_supprimer' => $nb_tags_supprimer );         }             $messages[] = $message;             $nb_erreur++;             $message['erreur'] = 1;             $message['message'] = __( "Erreur, aucun terms pour le post", TEXT_DOMAIN ) ;         {         else         }             }                 $messages[] = $message;                  }                     $nb_tags_supprimer++;                     $message['tags_supprimer'] = 1;                     $message['message'] = __( "Suppression du tag mais conservation de l'organisme ", TEXT_DOMAIN ) ;                 {                 else                 }                      $nb_supprimer++;                     $message['supprimer'] = 1;                     $message['message'] = __( "Suppression du tag et de l'organisme ", TEXT_DOMAIN );                      $this->_db->delete( $this->_db->posts, array( 'ID' => $post_id ) );                      // post organisme                      $this->_db->query( $this->_db->prepare( "DELETE FROM " . $this->_db->postmeta . " WHERE post_id = %s", $post_id ) );                       // meta datas                  {                 if( ! $terms_du_post ) // le post n'a plus aucun terms ( tag de la taxo taxo_tag )                 $terms_du_post = get_the_terms( $post_id, TAXO_TAG );                 // les terms du post                  $message = array( 'nom' => get_the_title( $post_id ), 'tag' => $slug_tag, 'message' => '', 'supprimer' => -1, 'tags_supprimer' => -1, 'erreur' => -1 );                 // message             {             foreach( $posts_id as $post_id )             // iterer a la recherche d'org orphelin                      wp_delete_term( $term_id, TAXO_TAG );             // supprimer le tag               $posts_id = get_objects_in_term( $term_id, TAXO_TAG );             // recuerer les orgs en rapport avec le tag              $term_id = $term->term_id;         {         if( $term )          $nb_erreur = 0;          $nb_tags_supprimer = 0;         $nb_supprimer = 0;         // les nb pour le message           $term = get_term_by( 'slug', $slug_tag, TAXO_TAG );         // recuperer l'id du term coorespondant au tag      {     public function supprimer_cpts( $slug_tag )     // supprimer      }         var_dump( $this->_db->last_query );     {     public function debug()    // utils      }         return $tags_formater;          }             $tags_formater = $tags_string;             $tags_string = substr( $tags_string, 0, -1 );             }                 $tags_string .= implode( ',', $tag_formater ) . ';' ;              {             foreach( $tags_formater as $tag_formater )             $tags_string = '';             // appartenance         {         if( $toString )          }             $tag_formater = array( 'tag_id' => $tag_id, 'tag_name' => $tag_name, 'tag_slug' => $tag_slug );              $tag_slug = ( array_key_exists( 'tag_slug', $tag ) ) ? $tag['tag_slug'] : false;             $tag_name = ( array_key_exists( 'tag_name', $tag ) ) ? $tag['tag_name'] : false;             $tag_id = ( array_key_exists( 'tag_id', $tag ) ) ? $tag['tag_id'] : false;         {         foreach( $tags as $tag )          $tags_formater = array();         // formater en tableau     {     public function formater_tags( $tags, $toString = false ) ad     �     g   �  �  �  n  J  $      �  �  �  �  �  �  h  Z      �  �  �  �  �  �  �  �  �      �  �  �  �  �  c  .    �  �  |    �
  �
  [
  #
  �	  �	  �  �  �  �  �  �  �  �  �  �  z  ]    �  �  �  �  �  �  �  �  z  @  ?      �  Z  P  	  �  �  �  �  �  d  E  ;  �  �  �  �  �  �  �  �  y  r  J       �  �  \  �  �  �                               *      * @param string $certification_active la certification qui est active ds le filtre ( on ne recupere que les cpt issut de celle la )      * @param string $ordre_trie ASC ou DESC      * @param string $order_by un nom de champ sur lequelle trier le resultat      * @param string $tag le nom du tag a utiliser ex charte_etic      *      * Recupere les posts_ids des cpt cpt      * Ne recupere pas l'id d'un cpt !!      *      * Recupere la liste des ids des custom post type cpt     /**      }         return $post_cpts;           }             $post_cpts[] = new $nom_class_api( $post_type, $id, 'localisation' );         {         foreach( $ids as $id )         $post_cpts = array();         $nom_class_api = ucfirst( $post_type ) . 'API'; // ex: OrganismeAPI          }             $ids = array( $post_id );         {         else // adresse unique ( ex afficahge de l'adresse d'un cpt );         }             $ids = $this->recuperer_posts_ids_cpt( $slug_tag, $post_type, 'post_title', 'ASC', 'string', $certification_active );             // recuperer une liste ( ex la map des cpt )         {         if( $post_id == false )          $post_id = ( $post_id == -1 ) ? false : $post_id;         // les js renvoient du -1 plutot que undefined ou false //FIXME bonne ou mvs idee ?!     {     public function recuperer_cpt_localisations( $slug_tag, $post_type, $post_id=false, $odre_trie = 'ASC', $certification_active = 'toute' ) // TODO refacto plus generic -> recupere cpt ( $post_type )      }          return $cpts;          }             $cpts[] = new $nom_class_api( $post_type, $id );             $nom_class_api = ucfirst( $post_type ) . 'API'; // ex: OrganismeAPI             $cpts = array();         {         if( $id )          //$this->debug();          }             // notify         {         else         }                 . "ORDER BY meta_value ASC", PREFIX_META . $nom_champ, $valeur_rechercher ) ); // TODO le PREFIX_META filtre deja les post type , ajouter quand mm une jointure pour filtre sur post_type explicitement ?                 . "AND meta_value = '%s' "                 . "WHERE meta_key = '%s' "                 . "FROM  " . $this->_db->postmeta . " "             $id = $this->_db->get_var( $this->_db->prepare( "SELECT DISTINCT post_id "             $nom_champ = 'nom_contact'; // fausse genericite // FIXME         {         else if( $nom_champ == 'nom_prenom_contact' ) // TODO concat nom prenom cas particulier nom_contact == nom prenom         }                 . "ORDER BY post_title ASC", $valeur_rechercher, $post_type ) );                 . "AND post_type = '%s' "                 . "WHERE post_title = '%s' "                 . "FROM  " . $this->_db->posts . " "             $id = $this->_db->get_var( $this->_db->prepare( "SELECT DISTINCT ID "         {         if( $nom_champ == 'post_title' )          $id = false;         $cpts = false;     {     public function recuperer_cpt_by_post_title_or_name_contact( $nom_champ, $valeur_rechercher, $post_type )      }         return $tags;          }             }                 $tags[] = $term->slug;             {             else             }                 $tags[Utils::get_id_tag( $term->slug )] = $term->slug;             {             if( $associatif )         {         foreach( $terms as $term )         $tags = array();         // transfo          $terms = get_terms( array( TAXO_TAG ), $args );          );             'cache_domain'  => 'core'             'search'        => '',              'offset'        => '',              'pad_counts'    => false,              'name__like'    => '',             'get'           => '',  