b0VIM 7.3      )D-T�  &  dendev                                  lt-devos                                /mnt/awt/dev-denis/organisme/wp-content/plugins/profil/src/admin/includes/Import.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �      ]         	      W         \   q            �         G   �         (   $                   D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ad  c  �     ]   �  �  �  �  �  }  `  ?  �  �  �  �  �  �  �  i  f  S  >        
  �  �  �  �  �    ~      �  �  �  �  �  &       �  �  �  �  o  i  h  2  ,       �
  �
  �
  }
  w
  v
  =
  7
  
  
  �	  �	  �	  ^	  ]	  ,	  �  �  �  E  ;  .  $  l  b  a  R  8  2  1    �  �  �  s  r  _  U  �  �  �  �  �  �  �  �  x  j  �  V  U  �  �  �  h    �  �  �  �      �  �  �           {         else         }             }                 $messages[] = array( 'message' => __( sprintf( 'Aucun %s de récupérer', $this->_post_type ), TEXT_DOMAIN ), 'type' => 'erreur' );             {             else             }                 update_option( DATE_IMPORT, $date_mise_a_jour );                 $date_mise_a_jour = $date_mise_a_jour->format( 'Y-m-d H:i:s' );                   $date_mise_a_jour = new DateTime('now',new DateTimeZone('Europe/London'));                 // conserver la date de mise a jour                  $messages = $this->_dbwp->ajouter_cpt( $cpt, $this->_post_type, $messages );                  $messages[] = array( 'message' => __( sprintf( 'le post type est : %s', $this->_post_type ) , TEXT_DOMAIN ), 'type' => 'debug' );                 $messages[] = array( 'message' => __( sprintf( 'le cpt : %s', $cpt_string ) , TEXT_DOMAIN ), 'type' => 'debug' );             {             if( $cpt )             // stocker en db wp              $cpt_string = print_r( $cpt, true );               }          }             $messages = $this->_dbwp->ajouter_cpt( $cpt, $this->_post_type, $messages );         {         if( $cpt )          update_option( 'mise_a_jour', $cpt );         $cpt = $this->_formater_import( $tmp_cpt, $this->_post_type );     {     public function mise_a_jour_cpt( $tmp_cpt )     // mise a jour      }         return $ids_cpts;         // fin          }             $messages[] = array( 'message' => __( sprintf( "Erreur: L'url ( %s ) d'acces au webservices est mauvaise", $this->_webservice_cpts  ), TEXT_DOMAIN ), 'type' => 'erreur' );         {         else         }             $messages[] = array( 'message' => __( sprintf( 'Il y a %s %s à importer',  count( $ids_cpts ), $nom_cpts ), TEXT_DOMAIN ), 'type' => 'info' );             // message              $ids_cpts = $rez->response->$nom_cpts;             $nom_cpts = $this->_post_type . 's';              $rez = json_decode( $rez_json );             $rez_json = file_get_contents( $this->_webservice_cpts );         {         if( $this->_verifier_url( $this->_webservice_cpts ) )          $ids_cpts = array();     {     public function recuperer_ids_cpts( &$messages ) //       }         return $this->_webservice_cpt;           $this->_webservice_cpt = URL_WEBSERVICE_CPTS . $id_cpt . '?oauth_token=' . $clee;          $clee = get_option( CLEE_IMPORT );     {     private function _url_detail_avec_clee( $id_cpt )      }         $this->_webservice_cpts = URL_WEBSERVICE_CPTS . 'listid?oauth_token=' . $clee;;          $clee = get_option( CLEE_IMPORT );     {     private function _url_avec_clee()      }         $this->_formatage_nom_db = array( 'id' => 'id_' . $this->_post_type, 'nom' => 'nom_' . $this->_post_type );         $this->_post_type = $post_type;           $this->_dbwp = Db::get_instance();          $this->_url_avec_clee();     {     public function __construct( $post_type ) // TODO parent et enfant profilImport pour la config ??        private $_post_type;     private $_formatage_nom_db;     private $_dbwp;     private $_webservice_cpt;     private $_webservice_cpts; { class Import  */  * @author   dendev <ddv@awt.be>  * @package  Options  * @category Admin  *  * Importe via la webservice les donnees cpts, tags, nomenclatures ds la db wp.  *  * Import ds wp des donnees de la db. /**    */  * @version  GIT: <http://magneto/stash/projects/WPPLO/repos/wp_plugin_cpt/browse>  * @author   dendev <ddv@awt.be>  * @package  WPPLO\Doc\Admin  *  * Permet de recuperer des cpts, tags, nomenclatures ds wp via le webservices.  *  * Liens entre wp et le webservice. /** <?php ad  �  �     D   �  �  �    �  �  �  �  T  >  �  �  �  e  G  �
  ^
  �	  �	  |	  5	  	  �  �  �  y  M  ;    �  �  �  �  �  �  P  F    	  �  �  �  ,  �  U  T      �  �  Z  @    �  �  �  �  q  @  2  (  '  &    �  �  �  �  �    t                                                                                                                                                                                                                                                                                                                                       ?> }?> }?>?> }     }         return $cpt;      ?> }     }         return $cpt;         print_r( $cpt );           }     ?> }     }         return $cpt;         print_r( $cpt );           }             }                 $cpt[$index] = $reseaux_sociaux;                 }                     }                         }                             $reseaux_sociaux[$nom] = $adresse;                         {                         else // url reseaux sociaux                         }                             $cpt['site_web_' . $nom_cpt] = $adresse;                         {                         if( strtolower( $nom ) == 'web' ) // url site web                     {                     if( $nom && $adresse && ! $lien_mort )                      $lien_mort = ( array_key_exists( 'lienMort', $tmp_url ) ) ? $tmp_url['lienMort'] : true;                     $adresse = ( array_key_exists( 'adresse', $tmp_url ) ) ? $tmp_url['adresse'] : false;                     $nom = ( array_key_exists( 'type', $tmp_url ) ) ? $tmp_url['type']['nom'] : false;                 {                 foreach( $tmp_cpt['urls'] as $tmp_url )                 $reseaux_sociaux = array();             {             if( is_array( $tmp_cpt['urls'] ) )         {         if( array_key_exists( 'urls', $tmp_cpt ) )         $cpt[$index] = false;         $index = 'reseaux_sociaux_' . $nom_cpt;         // reseaux sociaux          }             }                 $cpt['contact_contacts'] = $contacts;                 }                     $contacts[] = $contact;                     }                         }                             $contact['reseaux_sociaux'] = $reseaux_sociaux;                             }                                 }                                     $reseaux_sociaux[$nom] = $adresse;                                 {                                 if( $nom && $adresse && ! $lien_mort )                                 $lien_mort = ( array_key_exists( 'lienMort', $tmp_url ) ) ? $tmp_url['lienMort'] : true;                                 $adresse = ( array_key_exists( 'adresse', $tmp_url ) ) ? $tmp_url['adresse'] : false;                                 $nom = ( array_key_exists( 'type', $tmp_url ) ) ? $tmp_url['type']['nom'] : false;                             {                             foreach( $tmp_contact['urls'] as $tmp_url )                             $reseaux_sociaux = array();                         {                         if( is_array( $tmp_contact['urls'] ) )                     {                     if( array_key_exists( 'urls', $tmp_contact ) )                     $contact['reseaux_sociaux'] = false;                     // reseaux sociaux                     $contact['photo'] = ( array_key_exists( 'photo', $tmp_contact ) ) ? EMP_IMG_AWT . $tmp_contact['photo']['path'] : false;                     $contact['reseaux_sociaux'] = ( array_key_exists( 'reseaux_sociaux', $tmp_contact ) ) ? $tmp_contact['reseaux_sociaux'] : false;                     $contact['gsm'] = ( array_key_exists( 'gsm', $tmp_contact ) ) ? $tmp_contact['gsm'] : false;                     $contact['fax'] = ( array_key_exists( 'fax', $tmp_contact ) ) ? $tmp_contact['fax'] : false;                     $contact['telephone'] = ( array_key_exists( 'telephone', $tmp_contact ) ) ? $tmp_contact['telephone']['dial'] : false;                     $contact['prenom'] = ( array_key_exists( 'prenom', $tmp_contact ) ) ? $tmp_contact['prenom'] : false; ad  �  3     \   �  �  �  l  f  e  [  0  *      �  �  �  �  }  p  f  N  D  C  /  )  %  �  �  �  �  �  �  �    �  �  �    ~  0  �  �  �  �  �  �  �  �    m  J  �
  �
  �
  �
  `
  _
  A
  
  �	  �	  �	  R	  �  �  �  �  v  ;  1  �  �  �  �    �  3  �  �  �  �  t  j  i  Y  :    �  �  �  �  K  =  3  5  �  �  �  �  M  �  �                      // forme                     $entite_juridique['nom'] = ( array_key_exists( 'nom', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['nom'] : false;                     $entite_juridique['numero_tva'] = ( array_key_exists( 'numeroTVA', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['numeroTVA'] : false;                     $entite_juridique['numero_entreprise'] = ( array_key_exists( 'numeroEntreprise', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['numeroEntreprise'] : false;              $cpt[$index] = ( array_key_exists( 'logo', $tmp_cpt ) ) ? ( ( array_key_exists( 'path', $tmp_cpt['logo'] ) ) ? $tmp_cpt['logo']['path'        }             }                 $cpt[$index] = EMP_IMG_AWT . $tmp_cpt['logo']['path'];             {             if( array_key_exists( 'path', $tmp_cpt['logo'] ) )         {         if( array_key_exists( 'logo', $tmp_cpt ) )         $cpt[$index] = false;         $index = 'image_logo';         // logo          }             }                 $cpt[$index] = $presentation;                  );                     'de' => ( array_key_exists( 'de', $tmp_presentation ) ) ? $tmp_presentation['de'] : false                      'nl' => ( array_key_exists( 'nl', $tmp_presentation ) ) ? $tmp_presentation['nl'] : false,                     'en' => ( array_key_exists( 'en', $tmp_presentation ) ) ? $tmp_presentation['en'] : false,                 $presentation = array( 'fr' => ( array_key_exists( 'fr', $tmp_presentation ) ) ? $tmp_presentation['fr'] : false,                  $tmp_presentation = $tmp_cpt['presentation']['court'];             {             if( array_key_exists( 'court', $tmp_cpt['presentation'] ) )         {         if( array_key_exists( 'presentation', $tmp_cpt ) )         $cpt[$index] = false;         $index= 'description_' . $nom_cpt;         // description du cpt          $cpt[$index] = ( array_key_exists( 'dateModification', $tmp_cpt ) ) ? $tmp_cpt['dateModification'] : false;         $index = 'date_modification_' . $nom_cpt;         // date_modification_ cpt          $cpt[$index] = ( array_key_exists( 'dateCreation', $tmp_cpt ) ) ? $tmp_cpt['dateCreation'] : false;         $index = 'date_creation_' . $nom_cpt;         // date_creation_ cpt          $cpt[$index] = ( array_key_exists( 'nom', $tmp_cpt ) ) ? $tmp_cpt['nom'] : false;         $index = 'nom_' . $nom_cpt;         // nom cpt          $cpt[$index] = ( array_key_exists( 'id', $tmp_cpt ) ) ? $tmp_cpt['id'] : false;         $index = 'id_' . $nom_cpt;         // id cpt     {     private function _formater_import( $tmp_cpt, $nom_cpt )      }         return $cpt;           }             $cpt = $this->_formater_import( $cpt, $this->_post_type );             // formater ( recup les infos utils avec un index de nom formater              $cpt = $rez['response'][$this->_post_type];             // recupereation du cpt         {         if( is_array( $rez ) )         // recup les attributs de l'object sous forme d'un tableau, met le pointeur d'iteration au debut, demande la 1er cle          $rez = json_decode( $rez_json, true );         $rez_json = file_get_contents( $url );          $cpt = false;     {     private function _importer( $url )          }         return $ok;          }             $ok = $url;         {         else         }             $ok = false;         {         if( $url_headers[0] == 'HTTP/1.1 400 Bad Request' )          $url_headers = @get_headers( $url );          $ok = false;     {     private function _verifier_url( $url )     // --      }         return $items;          }             $messages[] = array( 'message' => __( 'Url paginée non valide', TEXT_DOMAIN ), 'type' => 'erreur' ); ad  �   �     G   �  r  \  
  �  �  �  p  B  �  �  �  J  �  l  �  �  k  M  0    �
  �
  M
  
  �	  2	  �  U  2      �  �  j  T  S  4  �  �  i  �  �  �  S    �  �  �  (    �  �  �  �  �  ]           �  �  �  b  T  /  �  �  �  �  �  �  t  j                $contact['nom'] = ( array_ke        }             }                 }                                                      $adresse = array();                 {                 foreach( $tmp_cpt['adresses'] as $tmp_adresse )                 $adresses = array();             {             if( is_array( $tmp_cpt['adresses'] ) )         {         if( array_key_exists( 'adresses', $tmp_cpt ) )         $cpt['adresse_adresses'] = false;         // adresses          }             $cpt['entites_juridiques'] = $entites_juridiques;             // ajout des infos entites juridique au infos cpts             }                 $entites_juridiques[] = $entite_juridique;                  }                     }                         }                             $entite_juridique['chiffres'] = $tmp_entite_juridique['chiffres'];                         {                         if( is_array( $tmp_entite_juridique['chiffres'] ) )                     {                     if( array_key_exists( 'chiffres', $tmp_entite_juridique ) )                     $entite_juridique['chiffres'] = false;                     // chiffres                      $entite_juridique['date_creation'] = ( array_key_exists( 'dateCreationOrganisme', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['dateCreationOrganisme'] : false;                     // date de creation juridique                      $entite_juridique['capital'] = ( array_key_exists( 'capital', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['capital'] : false;                     // capital                      }                         }                             $entite_juridique['forme'] = $forme;                             // ajouter la forme juridique aux infos juridique                              }                                 );                                     'de' => ( array_key_exists( 'de', $acronyme ) ) ? $acronyme['de'] : false                                     'nl' => ( array_key_exists( 'nl', $acronyme ) ) ? $acronyme['nl'] : false,                                     'en' => ( array_key_exists( 'en', $acronyme ) ) ? $acronyme['en'] : false,                                     'fr' => ( array_key_exists( 'fr', $acronyme ) ) ? $acronyme['fr'] : false,                                 $forme['acronyme'] = array(                                  $acronyme = $forme_juridique['acronyme'];                             {                             if( array_key_exists( 'acronyme', $forme_juridique ) )                             // acronyme                                                          }                                 );                                     'de' => ( array_key_exists( 'de', $intitule ) ) ? $intitule['de'] : false                                      'nl' => ( array_key_exists( 'nl', $intitule ) ) ? $intitule['nl'] : false,                                     'en' => ( array_key_exists( 'en', $intitule ) ) ? $intitule['en'] : false,                                     'fr' => ( array_key_exists( 'fr', $intitule ) ) ? $intitule['fr'] : false,                                 $forme['intitule'] = array(                                  $intitule = $forme_juridique['intitule'];                             {                             if( array_key_exists( 'intitule', $forme_juridique ) )                             $forme = array();                             // intitule                              $forme_juridique= $tmp_entite_juridique['formeJuridique'];                         {                         if( is_array( $tmp_entite_juridique['formeJuridique'] ) )                     {                     if( array_key_exists( 'formeJuridique', $tmp_entite_juridique ) )                     $entite_juridique['forme'] = false; ad    a        �  �  �  u  k  /  !  �  �  �  ]  �  
  ~  a  `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   // forme                     $entite_juridique['nom'] = ( array_key_exists( 'nom', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['nom'] : false;                     $entite_juridique['numero_tva'] = ( array_key_exists( 'numeroTVA', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['numeroTVA'] : false;                     $entite_juridique['numero_entreprise'] = ( array_key_exists( 'numeroEntreprise', $tmp_entite_juridique ) ) ? $tmp_entite_juridique['numeroEntreprise'] : false;                     $entite_juridique = array();                 {                 foreach( $tmp_cpt['entitesJuridiques'] as $tmp_entite_juridique )                 $entites_juridiques = array();             {             if( is_array( $tmp_cpt['entitesJuridiques'] ) )         {         if( array_key_exists( 'entitesJuridiques', $tmp_cpt ) )         $cpt['entites_juridiques'] = false;         // entites juridiques  ad  �  .        �  �  �  �  �  M  ?    �  �  �  �  .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            $contact['nom'] = ( array_key_exists( 'nom', $tmp_contact ) ) ? $tmp_contact['nom'] : false;                      $contact = array();                 {                 foreach( $tmp_cpt['contacts'] as $tmp_contact )                 $contacts = array();             {             if( is_array( $tmp_cpt['contacts'] ) )         {         if( array_key_exists( 'contacts', $tmp_cpt ) )         $cpt['contact_contacts'] = false;         // contacts  ad  3  �     (   �    �  !  �     �  r  /    �  �  Q  7  !     �
  �
  �
  E
  /
  �	  �	  j	  i	  	  �  �  a  C    �  �  �  o  C  1  #  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             }             $cpt['adresse_adresses'] = $adresses;             }                 }                     $adresses[] = $adresse;                     }                         }                             }                                 $adresse['longitude'] = $longitude;                                 $adresse['latitude'] = $latitude;                             {                             if( $latitude && $longitude )                              $longitude = ( array_key_exists( 1, $lat_long ) ) ? $lat_long[1] : false ;                             $latitude = ( array_key_exists( 0, $lat_long ) ) ? $lat_long[0] : false ;                              $lat_long = $tmp_adresse['position']['coordinates'];                         {                         if( array_key_exists( 'coordinates', $tmp_adresse['position'] ) )                     {                     if( array_key_exists( 'position', $tmp_adresse ) )                     $adresse['longitude'] = false;                     $adresse['latitude'] = false;                     // coordonnes geographique                      }                         }                             $adresse['pays'] = $tmp_adresse['pays']['localizedName'];                         {                         if( array_key_exists( 'localizedName', $tmp_adresse['pays'] ) )                     {                     if( array_key_exists( 'pays', $tmp_adresse ) )                     $adresse['pays'] = false;                     $adresse['localite'] = ( array_key_exists( 'localite', $tmp_adresse ) ) ? $tmp_adresse['localite'] : false;                     $adresse['code_postal'] = ( array_key_exists( 'codePostal', $tmp_adresse ) ) ? $tmp_adresse['codePostal'] : false;                     $adresse['numero'] = ( array_key_exists( 'numero', $tmp_adresse ) ) ? $tmp_adresse['numero'] : false;                     $adresse['rue'] = ( array_key_exists( 'rue', $tmp_adresse ) ) ? $tmp_adresse['rue'] : false;                     $adresse['principale'] = ( array_key_exists( 'principale', $tmp_adresse ) ) ? $tmp_adresse['principale'] : false;                     $adresse['type'] = ( array_key_exists( 'type', $tmp_adresse ) ) ? $tmp_adresse['type'] : false;                     $adresse['lieu'] = ( array_key_exists( 'lieu', $tmp_adresse ) ) ? $tmp_adresse['lieu'] : false; ad  j
  �
        �  �  �  �  �  f  4  *  �  �  �  �  �    �  k  j      �  }  +  �  �  �  �  )        �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    {         else         }             }                 $messages[] = array( 'message' => __( sprintf( 'Aucun %s de récupérer', $this->_post_type ), TEXT_DOMAIN ), 'type' => 'erreur' );             {             else             }                 update_option( DATE_IMPORT, $date_mise_a_jour );                 $date_mise_a_jour = $date_mise_a_jour->format( 'Y-m-d H:i:s' );                   $date_mise_a_jour = new DateTime('now',new DateTimeZone('Europe/London'));                 // conserver la date de mise a jour                  $messages = $this->_dbwp->ajouter_cpt( $cpt, $this->_post_type, $messages );                  $messages[] = array( 'message' => __( sprintf( 'le post type est : %s', $this->_post_type ) , TEXT_DOMAIN ), 'type' => 'debug' );                 $messages[] = array( 'message' => __( sprintf( 'le cpt : %s', $cpt_string ) , TEXT_DOMAIN ), 'type' => 'debug' );             {             if( $cpt )             // stocker en db wp              $cpt_string = print_r( $cpt, true );             $cpt = $this->_importer( $url_import );         {         if( $this->_verifier_url( $url_import ) )         $url_import = $this->_url_detail_avec_clee( $id_cpt );          $items = false;     {     public function importer_cpt( $id_cpt )     // importer 