b0VIM 7.3      �s�Sz   �  dendev                                  lt-devos                                /mnt/awt/dev-denis/agenda/wp-content/plugins/wp_plugin_agenda/src/commun/includes/cpts/CustomPostType.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �      k         ����U   l      ����o   �            0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ad  !   �     k   �  �  �  �  �  F  �  �  �  �  �  �  �  �  t  q  &  �  �  �  /  ,    �  �  �  �  �  �  �  �  L  F  6      �  �  ;  :  �
  �
  �
  �
  _
  �	  �	  �	  6	  5	  !	  �  b      �  �  �  �  �    1  �  �  }  v  :  2      �  �  �  u  k  6  ,      �  �  �  �  l  U  <  �  �  �  �  m  X  8  *              �  �  �  �  =  �  �  �  �                                    */      *      * @see http://codex.wordpress.org/Function_Reference/register_post_type      * callback appeler par la constructeur ( au travers d'un action wp )      * Utilise les informations de configuration pour la creation du cpt      *      * Creer un custom post type     /**      }         return $valeur;          }             }                 $valeur = true;             default:                 break;                 $valeur = $this->get_arg_config( 'slug' );             case 'post_type':                 break;                 $valeur = strtolower( $this->get_arg_config( 'nom' ) );             case 'slug':                 break;                 $valeur = 'test';             case 'nom':                 break;                 $valeur = 'post';             case 'capability_type':             {             switch( $nom )         {         else // renvoi une valeur par defaut adapter         }             $valeur = $this->_config[$nom];         {         if( array_key_exists( $nom, $this->_config ) )          // verifier si existe     {     public function get_arg_config( $nom )      */      * @return mixed la valeur de la configuration demander      *      * @param mixed[] $nom array associatif contenant les configurations a appliquer      *       * Si la config par defaut n'existe pas pour l'arg demander alors retrourne false.      * Si la configuration n'existe pas alors celle par defaut est appliquer.      * Retourne la valeur de la config demander via l'arguement.      *      * Recupere une des valeurs de la config.     /**      }         }             add_action( 'save_post', array( $nom_class_save, $nom_methode_save ) );             $nom_methode_save = strtolower( $this->get_arg_config( 'post_type' ) ) . '_save_callback';             $nom_class_save = ucfirst( $this->get_arg_config( 'post_type' ) ) . 'SAVE';             // save              add_action( 'load-post-new.php', array( $nom_class_render, $nom_methode_render ) );              add_action( 'load-post.php', array( $nom_class_render, $nom_methode_render ) );              $nom_methode_render = strtolower( $this->get_arg_config( 'post_type' ) ) . '_render_callback';             $nom_class_render = ucfirst( $this->get_arg_config( 'post_type' ) ) . 'RENDER';             // render         {          if( is_admin() )             // le render du cpt n'existe que pour l'interface admin           add_action( 'ajouter_supports', array( $this, 'ajouter_supports_callback' ), 10, 2 ); // supports d'edition: title, authors etc         add_action( 'init', array( $this, 'creer_cpt' )  );         // actions           $this->_config = $config;         // args     {     public function __construct( $config ) //TODO verifier l'args          private $_config; { abstract class CustomPostType //TODO abstract  */  * @author   dendev <ddv@awt.be>  * @package  Structure  * @category Organisme  *  * @param mixed[] $_config array associatif nom, valeur pour la configuration du cpt  *  * La personalisation se fait ds un enfant. CustomPostType n'est pas utiliser directement  * Et possibilite de rajouter des fonctionalites au custom post type  * Permet la creation d'un custom post type avec options de personlisation  *  * Crée un custom post type /**   */  * @author   dendev <ddv@awt.be>  * @package  Structure  * @category Organisme  *  * La personalisation se fait ds un enfant. CustomPostType n'est pas utiliser directement  * Et possibilite de rajouter des fonctionalites au custom post type  * Permet la creation d'un custom post type avec options de personlisation  *  * Crée un custom post type /** <?php ad  �
  �        �  j  '      �  �  �  �  �  �  H    P  ;  :    �  �  �  O    �  �  �  �  �  �  �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ?> }     }         wp_localize_script( 'sscpt-commun', 'sscpt', $js_vars );          }             );                 'sticky_count' => $sticky_count                 'sticky_text' => __( 'Sticky' ),                 'label_text' => __( 'Make this post sticky' ),                 'status_label_text' => __( 'Status' ),                 'post_type' => $screen->post_type,                 'screen' => 'edit',             $js_vars = array(                  : 0;                 ? $wpdb->get_var( $wpdb->prepare( "SELECT COUNT( 1 ) FROM $wpdb->posts WHERE post_type = %s AND post_status NOT IN ('trash', 'auto-draft') AND ID IN ($sticky_posts)", $screen->post_type ) )             $sticky_count = $sticky_posts             $sticky_posts = implode( ', ', array_map( 'absint', ( array ) get_option( 'sticky_posts' ) ) );              global $wpdb;         {         else          }              // Browsing custom posts              );                 'sticky_visibility_text' => __( 'Public, Sticky' )                 'label_text' => __( 'Stick this post to the front page' ),                 'checked_attribute' => checked( $is_sticky, true, false ), 