b0VIM 7.3      ġS�� �  dendev                                  lt-devos                                ~dendev/public_html/NeaLoca/wp-content/plugins/fmwp/fmwp.php                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 utf-8	 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �                  /            	   L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ad  s  �        �  �  �  �  �  >  ;  )    �  �  �  �  �  x  \  ?    �  �  �  �  w  l    �  �  M  �  �  �  C  �
  �
  5
  �	  �	  |	  (	  �  �  �  i        �  �  l  c    �  z  ,  +    �  �  }  t  #      �  �  _    �  B  �  �  |    �  h  g                                      	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/LocalisationSAVE.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/AccueilSAVE.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/CustomPostTypeSave.php';     // saves 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/ContactRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/ActiviteRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/AppartementRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/LocalisationRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/AccueilRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/AdminRENDER.php';     // renders 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/FmWpAdmin.php'; { if( is_admin() )   *----------------------------------------------------------------------------*/  * ADMIN /*----------------------------------------------------------------------------*  add_action( 'plugins_loaded', array( 'FmWpPublic', 'get_instance' ) ); // instancie le front  require_once plugin_dir_path( __FILE__ ) . 'src/public/includes/TestSHC.php'; require_once plugin_dir_path( __FILE__ ) . 'src/public/includes/ShortCode.php'; require_once plugin_dir_path( __FILE__ ) . 'src/public/FmWpPublic.php';  *----------------------------------------------------------------------------*/  * FRONT /*----------------------------------------------------------------------------*  add_action( 'plugins_loaded', array( 'FmWpCommun', 'get_instance' ) ); // instancie le commun  register_deactivation_hook( __FILE__, array( 'FmWpCommun', 'deactivate' ) ); register_activation_hook( __FILE__, array( 'FmWpCommun', 'activate' ) ); //activation et desactivation  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/psts/NealocaPST.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/psts/Posteur.php';  //posteur require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/ContactCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/ActiviteCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/AppartementCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/LocalisationCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/AccueilCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/CustomPostType.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/ApiCustomPostType.php'; /require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/AjaxHandler.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/Db.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/FmWpCommun.php'; require_once plugin_dir_path( __FILE__ ) . 'src/config.php';  *----------------------------------------------------------------------------*/  * COMMON  /*----------------------------------------------------------------------------*   */  * @license           GPL2   * Git Plugin URI:    https://github.com/nofh/fmwp.git  * Text Domain:       fmwp_lang  * Author:            dendev  * Version:           0.0.1  * Description:       Micro FrameWork  * Plugin URI:        @TODO  * Plugin Name:       NeaLoca   * @wordpress-plugin  *  * @author   dendev <ddv@awt.be>  * @package  Organisme  * @category Fmwp  *  * also follow WordPress Coding Standards and PHP best practices.  * A foundation off of which to build well-documented WordPress plugins that  *  * WordPress Micro FrameWork Plugin . /** <?php ad    ;     	   �  K  �  �  �  �  @  >  ;  :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ?> } 	add_action( 'plugins_loaded', array( 'FmWpAdmin', 'get_instance' ) );  	include_once plugin_dir_path( __FILE__ ) . 'src/admin/assets/vendors/simple_html_dom.php';     // vendors 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/ContactSAVE.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/ActiviteSAVE.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/AppartementSAVE.php'; ad  K       /   �  �  P  �  �  C  �  �  9  /  �  �  �  e    �  �  �  p  o      �
  }
  -
  �	  �	  �	  �	  �	  0	  '	  �  �  �  {  l    �  U  �  �  <  /  �  x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/LocalisationSAVE.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/AccueilSAVE.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/saves/CustomPostTypeSave.php';     // saves 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/ContactRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/ActiviteRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/AppartementRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/LocalisationRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/AccueilRENDER.php'; 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/includes/renders/AdminRENDER.php';     // renders 	include_once plugin_dir_path( __FILE__ ) . 'src/admin/FmWpAdmin.php'; { if( is_admin() )   *----------------------------------------------------------------------------*/  * ADMIN /*----------------------------------------------------------------------------*  add_action( 'plugins_loaded', array( 'FmWpPublic', 'get_instance' ) ); // instancie le front  require_once plugin_dir_path( __FILE__ ) . 'src/public/includes/TestSHC.php'; require_once plugin_dir_path( __FILE__ ) . 'src/public/includes/ShortCode.php'; require_once plugin_dir_path( __FILE__ ) . 'src/public/FmWpPublic.php';  *----------------------------------------------------------------------------*/  * FRONT /*----------------------------------------------------------------------------*  add_action( 'plugins_loaded', array( 'FmWpCommun', 'get_instance' ) ); // instancie le commun  register_deactivation_hook( __FILE__, array( 'FmWpCommun', 'deactivate' ) ); register_activation_hook( __FILE__, array( 'FmWpCommun', 'activate' ) ); //activation et desactivation  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/psts/NealocaPST.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/psts/Posteur.php';  //posteur require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/ContactCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/ActiviteCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/AppartementCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/LocalisationCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/AccueilCPT.php';  require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/CustomPostType.php'; require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/cpts/ApiCustomPostType.php'; //cpts require_once plugin_dir_path( __FILE__ ) . 'src/commun/includes/Utils.php'; 